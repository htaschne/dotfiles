library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity foo is
port(
    IN:  in  std_logic;
    OUT: out std_logic
);
end entity;

architecture arch of foo is
begin
    OUT <= (IN and OUT);
end architecture;
